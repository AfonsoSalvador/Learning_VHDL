library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity bin_counter is
   generic(N : integer := 32);
   
   port(
      clk      : in  std_logic;
      --reset    : in  std_logic;
      --enable   : in  std_logic;
      inc      : in std_logic; 
      dec      : in std_logic; 
      --max_tick : out std_logic;
      q        : out std_logic_vector(N-1 downto 0)
   );
end bin_counter;

architecture arch of bin_counter is
   signal r_reg  : unsigned(N-1 downto 0);
   signal r_next : unsigned(N-1 downto 0);
begin
   -- register
--   process(clk,reset)
--   begin
--      if (reset='1') then
--         r_reg <= (others=>'0');
--      elsif (clk'event and clk='1') then
--         if (enable='1') then
--            r_reg <= r_next;
--         end if;
--      end if;
--   end process;

process(clk)
   begin
      if (clk'event and clk='1') then
          r_reg <= r_next;
       end if;
   end process;
   
   
   -- next-state logic
   process(r_reg, inc, dec)
   begin
    if (inc='1') then 
        r_next <= r_reg + 1;
    
    elsif dec='1' then
        r_next <= r_reg - 1;
    else
        r_next <= r_reg;
    end if;
   
   end process;
   -- output logic
   q <= std_logic_vector(r_reg);
   --max_tick <= '1' when r_reg=(2**N - 1) else '0';
end arch;