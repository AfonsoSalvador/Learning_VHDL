library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity free_run_bin_counter is
   generic(N : integer := 15);
   --generic(N : integer := 8);
   port(
      clk      : in  std_logic;
      reset    : in  std_logic;
      enable   : in  std_logic;
      max_tick : out std_logic;
      q        : out std_logic_vector(N-1 downto 0)
   );
end free_run_bin_counter;

architecture arch of free_run_bin_counter is
   signal r_reg  : unsigned(N-1 downto 0); -- registrador 
   signal r_next : unsigned(N-1 downto 0); -- mudança de estado 
begin
   -- register
   process(clk,reset)
   begin
      if (reset='1') then
         r_reg <= (others=>'0');
      elsif (clk'event and clk='1') then -- se tiver um evento de clock e for uma borda de subida 
         if (enable='1') then
            r_reg <= r_next;
         end if;
      end if;
   end process;
   -- next-state logic
   r_next <= r_reg + 1; -- estado atual + 1 
   -- output logic
   q <= std_logic_vector(r_reg);
   max_tick <= '1' when r_reg=(2**N - 1) else '0'; -- só é um quando o registrador alcança o valor máximo 
end arch;